// Zuhair Shaikh and Brant Lan Li
// ADD Operation (ADD)
// ELEC374 - Digital Systems Engineering
// Department of Electrical and Computer Engineering
// Queen's University

module adder_4(
	input wire [3:0] rA, rB,
	input wire cIn,
	output wire [3:0] S,
	output wire cOut
	);
	
	wire [3:0] G;
	wire [3:0] P; 
	wire [3:0] C;
	
	assign G = rA ^ rB;
	assign P = rA & rB;
	assign C[0] = cIn;
	assign C[1]= G[0] | (P[0]&C[0]);
	assign C[2]= G[1] | (P[1]&G[0]) | P[1]&P[0]&C[0];
	assign C[3]= G[2] | (P[2]&G[1]) | P[2]&P[1]&G[0] | P[2]&P[1]&P[0]&C[0];
	assign cout = G[3] | (P[3]&G[2]) | P[3]&P[2]&G[1] | P[3]&P[2]&P[1]&G[0] | P[3]&P[2]&P[1]&P[0]&C[0];
	assign S[3:0] = P ^ C;
endmodule

module adder_16(
	input wire [15:0] rA, rB,
	input wire cIn,
	output wire [15:0] S,
	output wire cOut
	);
	
	wire cOutA;
	wire cOutB;
	wire cOutC;

	adder_4 adderA(.rA(rA[3:0]), .rB(rB[3:0]), .cIn(cIn), .S(S[3:0]), .cOut(cOutA));
	adder_4 adderB(.rA(rA[7:4]), .rB(rB[7:4]), .cIn(cOutA), .S(S[7:4]), .cOut(cOutB));				
	adder_4 adderC(.rA(rA[11:8]), .rB(rB[11:8]), .cIn(cOutB), .S(S[11:8]), .cOut(cOutC));
	adder_4 adderD(.rA(rA[15:12]), .rB(rB[15:12]), .cIn(cOutC), .S(S[15:12]), .cOut(cOut));
endmodule

module adder_32(
	input wire [31:0] rA, rB,
	input wire cIn,
	output wire [31:0] S,
	output wire cOut
	);
	
	wire cOutTemp;

	adder_16 adderA(.rA(rA[15:0]), .rB(rB[15:0]), .cIn(cIn), .S(S[15:0]), .cOut(cOutTemp));
	adder_16 adderB(.rA(rA[31:16]), .rB(rB[31:16]), .cIn(cOutTemp), .S(S[31:16]), .cOut(cOut));
endmodule